*** SPICE deck for cell flip_flop_MS{lay} from library D_flip_flop_MS
*** Created on Thu May 20, 2021 13:41:11
*** Last revised on Thu May 20, 2021 14:37:05
*** Written on Sun Oct 03, 2021 10:48:27 by Electric VLSI Design System,
*version 9.00
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: flip_flop_MS{lay}
Mnmos@0 net@5 D gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U PD=6U
Mnmos@1 net@15 CLK net@5 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U PD=9.5U
Mnmos@2 net@38 CLK gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U PD=6U
Mnmos@3 net@34 net@49 net@38 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U
+PD=9.5U
Mnmos@4 net@49 D gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=10.125P PS=32.7U
+PD=13.5U
Mnmos@5 net@70 net@15 gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U
+PD=6U
Mnmos@6 net@66 net@78 net@70 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U
+PD=9.5U
Mnmos@7 net@82 net@66 gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U
+PD=6U
Mnmos@8 net@78 net@34 net@82 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U
+PD=9.5U
Mnmos@9 net@230 net@66 gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U
+PD=6U
Mnmos@10 net@199 net@185 net@230 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U
+PD=9.5U
Mnmos@11 net@237 net@185 gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U
+PD=6U
Mnmos@12 net@211 net@78 net@237 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U
+PD=9.5U
Mnmos@13 net@246 net@199 gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U
+PD=6U
Mnmos@14 Q Qbar net@246 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U PD=9.5U
Mnmos@15 net@253 Q gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=4.5P PS=32.7U PD=6U
Mnmos@16 Qbar net@211 net@253 gnd NMOS L=0.6U W=3U AS=4.5P AD=8.25P PS=6U
+PD=9.5U
Mnmos@17 net@185 CLK gnd gnd NMOS L=0.6U W=3U AS=22.95P AD=10.125P PS=32.7U
+PD=13.5U
Mpmos@0 net@15 D vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P PS=28.833U
+PD=9.5U
Mpmos@1 vdd CLK net@15 vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U
+PD=28.833U
Mpmos@2 net@34 CLK vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P PS=28.833U
+PD=9.5U
Mpmos@3 vdd net@49 net@34 vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U
+PD=28.833U
Mpmos@4 net@49 D vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=10.125P PS=28.833U
+PD=13.5U
Mpmos@5 net@66 net@15 vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P PS=28.833U
+PD=9.5U
Mpmos@6 vdd net@78 net@66 vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U
+PD=28.833U
Mpmos@7 net@78 net@66 vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P PS=28.833U
+PD=9.5U
Mpmos@8 vdd net@34 net@78 vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U
+PD=28.833U
Mpmos@9 net@199 net@66 vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P PS=28.833U
+PD=9.5U
Mpmos@10 vdd net@185 net@199 vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U
+PD=28.833U
Mpmos@11 net@211 net@185 vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P
+PS=28.833U PD=9.5U
Mpmos@12 vdd net@78 net@211 vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U
+PD=28.833U
Mpmos@13 Q net@199 vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P PS=28.833U
+PD=9.5U
Mpmos@14 vdd Qbar Q vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U PD=28.833U
Mpmos@15 Qbar Q vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=8.25P PS=28.833U PD=9.5U
Mpmos@16 vdd net@211 Qbar vdd PMOS L=0.6U W=6U AS=8.25P AD=22.5P PS=9.5U
+PD=28.833U
Mpmos@17 net@185 CLK vdd vdd PMOS L=0.6U W=6U AS=22.5P AD=10.125P PS=28.833U
+PD=13.5U

* Spice Code nodes in cell cell 'flip_flop_MS{lay}'
vdd vdd 0 DC 5
vin D 0 pulse 0 5 2m 1n 1n 8m 16m
vin2 CLK 0 pulse 0 5 1m 1n 1n 4m 8m
.tran 24m
.include C5_models.txt
.END
