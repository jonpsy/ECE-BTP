*** SPICE deck for cell GDI{lay} from library GDI
*** Created on Tue Sep 21, 2021 15:25:54
*** Last revised on Tue Sep 21, 2021 16:28:24
*** Written on Tue Sep 21, 2021 16:29:10 by Electric VLSI Design System,
*version 9.00
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2
*** WARNING: no power connection for P-transistor wells in cell
*'GDI:GDI{lay}'

*** TOP LEVEL CELL: GDI:GDI{lay}
Mnmos@1 D G gnd gnd NMOS L=0.6U W=3U AS=20.25P AD=10.125P PS=31.5U PD=13.5U
Mpmos@1 D G P vdd PMOS L=0.6U W=6U AS=22.5P AD=10.125P PS=31.5U PD=13.5U

* Spice Code nodes in cell cell 'GDI:GDI{lay}'
vin G 0 pulse 0 5 0 1n 1n 8m 16m
vin2 P 0 pulse 0 5 0 1n 1n 4m 8m
.tran 16m
.include C5_models.txt
.END
