*** SPICE deck for cell GDI-DFF{lay} from library GDI
*** Created on Tue Sep 28, 2021 12:42:43
*** Last revised on Thu Sep 30, 2021 16:43:43
*** Written on Thu Sep 30, 2021 17:05:27 by Electric VLSI Design System,
*version 9.00
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: GDI-DFF{lay}
Mnmos@0 net@29 net@177 gnd gnd NMOS L=0.6U W=3U AS=43.65P AD=10.125P PS=53.7U
+PD=13.5U
Mnmos@8 net@168 net@215 gnd gnd NMOS L=0.6U W=3U AS=43.65P AD=10.125P
+PS=53.7U PD=13.5U
Mnmos@9 net@177 CLK net@168 gnd NMOS L=0.6U W=3U AS=10.125P AD=10.125P
+PS=13.5U PD=13.5U
Mnmos@10 net@215 CLK net@29 gnd NMOS L=0.6U W=3U AS=10.125P AD=10.125P
+PS=13.5U PD=13.5U
Mnmos@11 net@376 CLK Q gnd NMOS L=0.6U W=3U AS=9P AD=10.125P PS=12.5U
+PD=13.5U
Mnmos@12 Q_BAR net@376 gnd gnd NMOS L=0.6U W=3U AS=43.65P AD=9P PS=53.7U
+PD=12.5U
Mnmos@13 net@420 CLK Q_BAR gnd NMOS L=0.6U W=3U AS=9P AD=10.125P PS=12.5U
+PD=13.5U
Mnmos@14 Q net@420 gnd gnd NMOS L=0.6U W=3U AS=43.65P AD=9P PS=53.7U PD=12.5U
Mpmos@0 net@29 net@177 vdd vdd PMOS L=0.6U W=6U AS=51.3P AD=10.125P PS=60.3U
+PD=13.5U
Mpmos@9 net@177 CLK D vdd PMOS L=0.6U W=6U AS=13.5P AD=10.125P PS=16.5U
+PD=13.5U
Mpmos@10 net@215 CLK D_BAR vdd PMOS L=0.6U W=6U AS=13.5P AD=10.125P PS=16.5U
+PD=13.5U
Mpmos@11 net@376 CLK net@168 vdd PMOS L=0.6U W=6U AS=10.125P AD=10.125P
+PS=13.5U PD=13.5U
Mpmos@12 Q_BAR net@376 vdd vdd PMOS L=0.6U W=6U AS=51.3P AD=9P PS=60.3U
+PD=12.5U
Mpmos@13 net@420 CLK net@29 vdd PMOS L=0.6U W=6U AS=10.125P AD=10.125P
+PS=13.5U PD=13.5U
Mpmos@14 Q net@420 vdd vdd PMOS L=0.6U W=6U AS=51.3P AD=9P PS=60.3U PD=12.5U
Mpmos@15 net@168 net@215 vdd vdd PMOS L=0.6U W=6U AS=51.3P AD=10.125P
+PS=60.3U PD=13.5U

* Spice Code nodes in cell cell 'GDI-DFF{lay}'
vdd vdd 0 DC 5
vin D 0 pulse 0 5 2m 1n 1n 8m 16m
vin2 D_BAR 0 pulse 5 0 2m 1n 1n 8m 16m
vin3 CLK 0 pulse 0 5 1m 1n 1n 4m 8m
.tran 24m
.include C5_models.txt
.END
